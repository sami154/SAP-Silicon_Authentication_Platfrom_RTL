`timescale 1ns/1ps
module tb_PUF();
localparam    CHALLENGE_SIZE = 32,
              RESPONSE_SIZE = 256,
              HELPER_DATA_SIZE = 96;

	reg [CHALLENGE_SIZE-1:0] CHALLENGE;
	reg CLK;
	reg RST;
	reg INPUT_READY;
	reg [0:HELPER_DATA_SIZE-1] HELPER_DATA;
	wire [RESPONSE_SIZE-1:0] PUF_RESPONSE;
	wire DONE;



always #10 CLK = ~CLK;

initial begin

	CLK = 0;
	RST = 1;
	#20;
	RST = 0;
	INPUT_READY = 0;
	HELPER_DATA = 0;
	CHALLENGE = 'd0;
	#20;
	CHALLENGE = 'd1;
	HELPER_DATA = 96'b000001111001011010110101010110011111111101000010011101101000111110100101111100011111101111000101;
//	HELPER_DATA = 96'b0;
	#20;
	INPUT_READY = 1;
	#20;
	INPUT_READY = 0;
	wait(DONE == 1);
	$display("PUF PUF_RESPONSE 1: %h", PUF_RESPONSE);
	#300;
	CHALLENGE = 'd3;
//	HELPER_DATA = 96'b000001111001011010110101010110011111111101000010011101101000111110100101111100011111101111000101;
	HELPER_DATA = 96'b0;
	#20;
	INPUT_READY = 1;
	#20;
	INPUT_READY = 0;
	#500;
//	$display("PUF PUF_RESPONSE 2: %h", PUF_RESPONSE);

	


end

	wrapper_puf #(
				.CHALLENGE_SIZE(CHALLENGE_SIZE),
	            .RESPONSE_SIZE(RESPONSE_SIZE),
                .HELPER_DATA_SIZE(HELPER_DATA_SIZE)
	
	) WR_PUF ( 
				.CHALLENGE(CHALLENGE),
				.CLK(CLK),
				.RST(RST),
				.INPUT_READY(INPUT_READY),
				.HELPER_DATA(HELPER_DATA),
				.PUF_RESPONSE(PUF_RESPONSE),
				.DONE(DONE)
	
	);


endmodule